module comparador(
    input  logic [6:0] data_paridad, 
    input  logic [6:0] comparacion
);
endmodule

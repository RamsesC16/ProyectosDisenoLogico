module comparador(
    logic [6:0] data_paridad, 
    logic [6:0] comparacion,

)
endmodule